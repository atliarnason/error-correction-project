-- -----------------------------------------------------------------------------
--
--  Title      :  Testbench for Hamming SEC-DED decoder
--             :
--  Purpose    :  Non-exhaustive test of decoder
--             :
-- -----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_textio.all;

use work.Util.all;

entity HammingDecoderTb is
end entity;

architecture TestBench of HammingDecoderTb is 

    component HammingDecoder is 
        port(
            x_encoded:  in  std_logic_vector(7 downto 0);
            x:          out std_logic_vector(3 downto 0);
            corrected:  out std_logic;
error:      out std_logic
        );
    end component;

    signal encoded:  std_logic_vector(7 downto 0) := "00000000";
    signal decoded, expected: std_logic_vector(3 downto 0) := "0000";
    signal corrected, error: std_logic := '0';

begin

    dut: HammingDecoder 
        port map(
            x_encoded => encoded, 
            x => decoded,
            corrected => corrected,
            error => error
        );

    


    process
        constant period: time := 200 ns;
    begin
       

        -- Testing will test 3 category of cases: no noise, 1 error and 2 errors
        -- Test-cases can be generated with little effort using Python


        -- Testing messages with no artificial errors.
        -- Shows what encoded message is being input, and then complains if there is an error.
        
        -- ######################################### --
        -- ####### AUTOGENERATED WITH PYTHON ####### --
        -- ######################################### --

        encoded <= "00000000";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "0000"))
		    report("Test failed for " & "00000000" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "10000111";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "0001"))
		    report("Test failed for " & "10000111" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "10011001";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "0010"))
		    report("Test failed for " & "10011001" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "00011110";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "0011"))
		    report("Test failed for " & "11110000" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "10101010";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "0100"))
		    report("Test failed for " & "10101010" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "00101101";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "0101"))
		    report("Test failed for " & "10110100" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "00110011";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "0110"))
		    report("Test failed for " & "11001100" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "10110100";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "0111"))
		    report("Test failed for " & "10110100" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "01001011";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "1000"))
		    report("Test failed for " & "10010110" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "11001100";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "1001"))
		    report("Test failed for " & "11001100" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "11010010";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "1010"))
		    report("Test failed for " & "11010010" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "01010101";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "1011"))
		    report("Test failed for " & "10101010" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "11100001";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "1100"))
		    report("Test failed for " & "11100001" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "01100110";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "1101"))
		    report("Test failed for " & "11001100" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "01111000";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "1110"))
		    report("Test failed for " & "11110000" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));

	    encoded <= "11111111";
	    wait for period;
	    report( "Encoded message is " & to_string(encoded));
	    assert ((corrected = '0') and (error = '0') and (decoded = "1111"))
		    report("Test failed for " & "11111111" & " | Corrected or Error are wrong: " & to_string(corrected) & to_string(error));


        -- Add artificial noise. A random noise mask will be xor'ed with each encoded message.
        -- This mask will have 1 hi bit, resulting in 1 error occurring. (exhaustive testing of 
        -- this would require 128 test cases.)









        wait; -- indefinitely suspend process
    end process;

end architecture;
